`timescale 1ns/100ps


//CALCULATES THE ADDITIONAL J,BEQ,BNE SHIFT VALUE
//IN THIS MODULE 
//J,BEQ,BNE  ADDER IS CALLED HERE
//BY CHECKING WITH ZERO THE LAST SHIFTING VALUE OUTPUTS HERE.
module add(SHIFTS,J,BEQ,BNE,ZERO, PC_INC);

    //INITILIZE INPUTS
    input J,BEQ,BNE,ZERO;
    input [7:0] SHIFTS;
    input [31:0] PC;
    //INITILIZE OUTPUT
    output reg [31:0] PC_INC=32'b0;

    reg OUT1,OUT2,OUT3,OUT4;//SIGNALS
    reg [31:0] CHECK;//1 VALUE  IF SHIFT POSSIBLE ELSE 0
    reg [31:0] ADD;  
    wire [31:0] CAL_SHIFTS;//STORES OFFSET CALCULATED BY shift_adder  BELOW
   
    
    always@(*)
    begin
        
        // CHECK IF SHOULD SHIFTED
        OUT1=BEQ &&  ZERO; // IF BEQ
        OUT2=BNE && ~ZERO;//BNE
        OUT3=OUT2||OUT1;
        OUT4=OUT3||J;
        CHECK=$signed(OUT4);
        
        //REAL VALUE TO SHIFT AFTER CHECKING FOR ZERO
        //AND THE 0 OR 1 VALUE WITH PRE CALCULATED CAL_SHIFTS
        ADD=CHECK & CAL_SHIFTS;
        //MAKE ADD TO 32 BITS
        PC_INC= ADD;


    end
    
    //ADDITIONAL J,BEQ,BNE OFFSET VALUE IS CALCULATED HERE
    //THIS ADDER WORKS  AFTER INSTRUCTION MEMORY READ AND PARALLEL TO REG READ .
    //RETURNS OFFSET WITH #2 DELAY
    //MODULE IS AT two_adders.v
    //CAL_SHIFT STORES OFFSET
    shift_adder shifts(SHIFTS,CAL_SHIFTS);
endmodule